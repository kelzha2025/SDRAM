/////////////////////////////////////////////////////////////////
////        This is the package file.                        ////
////                                                         ////
////                                                         ////
////     Created By: Manasa Gurrala                          ////
////                 Venkata Naveen Reddy Yalla              ////
////                 Karthik Rudraraju                       ////
////                                                         ////
/////////////////////////////////////////////////////////////////

package sdrctrl_package;
import uvm_pkg::*;
import tb_classes_pkg::*;
`include "uvm_macros.svh"


endpackage : sdrctrl_package
