/////////////////////////////////////////////////////////////////
////        This is the package file.                        ////
////                                                         ////
////                                                         ////
////     Created By: Manasa Gurrala                          ////
////                 Venkata Naveen Reddy Yalla              ////
////                 Karthik Rudraraju                       ////
////                                                         ////
/////////////////////////////////////////////////////////////////

package sdrctrl_package;
import uvm_pkg::*;

`include "uvm_macros.svh"
// Core transaction and agent components
`include "sdr_seq_item.svh"
`include "sdr_sequence.svh"
`include "sdr_sequencer.svh"
`include "sdr_driver.svh"
`include "sdr_monitor.svh"
`include "sdr_agent.svh"
`include "cov_adapter.svh"

// Legacy/testbench utilities
`include "coverage.svh"
`include "stimulus_tester.svh"
`include "stimulus_values.svh"
`include "scoreboard.svh"
`include "env.svh"
`include "test.svh"


endpackage : sdrctrl_package
