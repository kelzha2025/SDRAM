package coverage_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "coverage.svh"
endpackage : coverage_pkg
