package tb_classes_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  import coverage_pkg::*;
  `include "sdr_seq_item.svh"
  `include "sdr_sequence.svh"
  `include "sdr_sequencer.svh"
  `include "sdr_driver.svh"
  `include "sdr_monitor.svh"
  `include "sdr_agent.svh"
  `include "cov_adapter.svh"
  `include "scoreboard.svh"
  `include "stimulus_tester.svh"
  `include "stimulus_values.svh"
  `include "env.svh"
  `include "test.svh"
endpackage : tb_classes_pkg
